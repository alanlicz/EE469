// a shifter,  by deflaut take 32 input width, output 32 output width
module shifterP #(parameter WIDTH = 32) (
	input logic		[WIDTH-1:0]	value,
	input logic					direction, // 0: left, 1: right
	input	logic		[5:0]		distance,  //shamt
	output logic	[WIDTH-1:0]	result
	);
	
	always_comb begin
		if (direction == 0)
			result = value << distance;
		else
			result = value >> distance;
	end
endmodule 